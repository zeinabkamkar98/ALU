`timescale 1ns / 1ps

module ieee_tes(
    );


endmodule
